magic
tech ihp-sg13g2
timestamp 1746729020
<< poly >>
rect 0 786 50 793
rect 0 770 7 786
rect 43 770 50 786
rect 0 750 50 770
rect 0 -20 50 0
rect 0 -36 7 -20
rect 43 -36 50 -20
rect 0 -43 50 -36
<< polycont >>
rect 7 770 43 786
rect 7 -36 43 -20
<< xpolyres >>
rect 0 0 50 750
<< metal1 >>
rect 2 786 48 791
rect 2 770 7 786
rect 43 770 48 786
rect 2 765 48 770
rect 2 -20 48 -15
rect 2 -36 7 -20
rect 43 -36 48 -20
rect 2 -41 48 -36
<< labels >>
flabel comment s 25 375 25 375 0 FreeSans 100 90 0 0 rpnd r=22493.913
<< end >>
