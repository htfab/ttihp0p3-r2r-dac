magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746729020
<< metal1 >>
rect 18935 27306 19035 27315
rect 18935 27229 18936 27306
rect 19034 27229 19035 27306
rect 18935 27221 19035 27229
rect 20111 27306 20211 27315
rect 20111 27229 20112 27306
rect 20210 27229 20211 27306
rect 20111 27221 20211 27229
rect 21287 27306 21387 27315
rect 21287 27229 21288 27306
rect 21386 27229 21387 27306
rect 21287 27221 21387 27229
rect 22463 27306 22563 27315
rect 22463 27229 22464 27306
rect 22562 27229 22563 27306
rect 22463 27221 22563 27229
rect 23999 26724 24439 26733
rect 23999 26622 24000 26724
rect 23247 26394 24000 26622
rect 23999 26284 24000 26394
rect 24438 26284 24439 26724
rect 23999 26275 24439 26284
rect 18601 25815 18781 25823
rect 18543 25814 18839 25815
rect 18347 25720 18447 25729
rect 18347 25643 18348 25720
rect 18446 25643 18447 25720
rect 18347 25635 18447 25643
rect 18543 25636 18602 25814
rect 18780 25636 18839 25814
rect 18543 25635 18839 25636
rect 19523 25720 19623 25729
rect 19523 25643 19524 25720
rect 19622 25643 19623 25720
rect 19523 25635 19623 25643
rect 20699 25720 20799 25729
rect 20699 25643 20700 25720
rect 20798 25643 20799 25720
rect 20699 25635 20799 25643
rect 21875 25720 21975 25729
rect 21875 25643 21876 25720
rect 21974 25643 21975 25720
rect 21875 25635 21975 25643
rect 18601 25627 18781 25635
<< via1 >>
rect 18936 27229 19034 27306
rect 20112 27229 20210 27306
rect 21288 27229 21386 27306
rect 22464 27229 22562 27306
rect 24000 26284 24438 26724
rect 18348 25643 18446 25720
rect 18602 25636 18780 25814
rect 19524 25643 19622 25720
rect 20700 25643 20798 25720
rect 21876 25643 21974 25720
<< metal2 >>
rect 18358 30266 18436 30274
rect 18348 30186 18357 30266
rect 18437 30186 18446 30266
rect 18358 30178 18436 30186
rect 18367 25720 18427 30178
rect 18946 29868 19024 29876
rect 18936 29788 18945 29868
rect 19025 29788 19034 29868
rect 18946 29780 19024 29788
rect 18955 27306 19015 29780
rect 19534 29466 19612 29474
rect 19524 29386 19533 29466
rect 19613 29386 19622 29466
rect 19534 29378 19612 29386
rect 18927 27229 18936 27306
rect 19034 27229 19043 27306
rect 18601 25814 18781 25815
rect 18339 25643 18348 25720
rect 18446 25643 18455 25720
rect 18593 25636 18602 25814
rect 18780 25636 18789 25814
rect 19543 25720 19603 29378
rect 20122 29066 20200 29074
rect 20112 28986 20121 29066
rect 20201 28986 20210 29066
rect 20122 28978 20200 28986
rect 20131 27306 20191 28978
rect 20710 28666 20788 28674
rect 20700 28586 20709 28666
rect 20789 28586 20798 28666
rect 20710 28578 20788 28586
rect 20103 27229 20112 27306
rect 20210 27229 20219 27306
rect 20719 25720 20779 28578
rect 21298 28266 21376 28274
rect 21288 28186 21297 28266
rect 21377 28186 21386 28266
rect 21298 28178 21376 28186
rect 21307 27306 21367 28178
rect 21886 27866 21964 27874
rect 21876 27786 21885 27866
rect 21965 27786 21974 27866
rect 21886 27778 21964 27786
rect 21279 27229 21288 27306
rect 21386 27229 21395 27306
rect 21895 25720 21955 27778
rect 22474 27466 22552 27474
rect 22464 27386 22473 27466
rect 22553 27386 22562 27466
rect 22473 27306 22553 27386
rect 22455 27229 22464 27306
rect 22562 27229 22571 27306
rect 24000 26724 24440 26733
rect 23991 26284 24000 26724
rect 24440 26284 24447 26724
rect 24000 26275 24440 26284
rect 19515 25643 19524 25720
rect 19622 25643 19631 25720
rect 20691 25643 20700 25720
rect 20798 25643 20807 25720
rect 21867 25643 21876 25720
rect 21974 25643 21983 25720
rect 18601 24776 18781 25636
rect 18592 24596 18601 24776
rect 18781 24596 18790 24776
rect 18601 24589 18781 24596
<< via2 >>
rect 18357 30186 18437 30266
rect 18945 29788 19025 29868
rect 19533 29386 19613 29466
rect 20121 28986 20201 29066
rect 20709 28586 20789 28666
rect 21297 28186 21377 28266
rect 21885 27786 21965 27866
rect 22473 27386 22553 27466
rect 24000 26284 24438 26724
rect 24438 26284 24440 26724
rect 18601 24596 18781 24776
<< metal3 >>
rect 18357 30266 18437 30275
rect 30500 30256 30556 30263
rect 18437 30196 30498 30256
rect 30558 30196 30567 30256
rect 30500 30189 30556 30196
rect 18357 30177 18437 30186
rect 18945 29868 19025 29877
rect 31266 29858 31326 29867
rect 19025 29798 31266 29858
rect 31266 29789 31326 29798
rect 18945 29779 19025 29788
rect 19533 29466 19613 29475
rect 32034 29456 32094 29465
rect 19613 29396 32034 29456
rect 32034 29387 32094 29396
rect 19533 29377 19613 29386
rect 20121 29066 20201 29075
rect 32802 29056 32862 29065
rect 20201 28996 32802 29056
rect 32802 28987 32862 28996
rect 20121 28977 20201 28986
rect 20709 28666 20789 28675
rect 33570 28656 33630 28665
rect 20789 28596 33570 28656
rect 33570 28587 33630 28596
rect 20709 28577 20789 28586
rect 21297 28266 21377 28275
rect 34338 28256 34398 28265
rect 21377 28196 34338 28256
rect 34338 28187 34398 28196
rect 21297 28177 21377 28186
rect 21885 27866 21965 27875
rect 35106 27856 35166 27865
rect 21965 27796 35106 27856
rect 35106 27787 35166 27796
rect 21885 27777 21965 27786
rect 22473 27466 22553 27475
rect 35874 27456 35934 27465
rect 22553 27396 35874 27456
rect 35874 27387 35934 27396
rect 22473 27377 22553 27386
rect 24000 26724 24440 26733
rect 23991 26284 24000 26724
rect 24440 26284 24449 26724
rect 24000 26275 24440 26284
rect 620 24776 800 24785
rect 18601 24776 18781 24785
rect 800 24596 18601 24776
rect 620 24587 800 24596
rect 18601 24587 18781 24596
<< via3 >>
rect 30498 30196 30558 30256
rect 31266 29798 31326 29858
rect 32034 29396 32094 29456
rect 32802 28996 32862 29056
rect 33570 28596 33630 28656
rect 34338 28196 34398 28256
rect 35106 27796 35166 27856
rect 35874 27396 35934 27456
rect 24000 26284 24440 26724
rect 620 24596 800 24776
<< metal4 >>
rect 5913 30797 5922 30857
rect 5982 30797 5991 30857
rect 5922 30596 5982 30797
rect 6681 30796 6690 30856
rect 6750 30796 6759 30856
rect 7449 30796 7458 30856
rect 7518 30796 7527 30856
rect 8217 30796 8226 30856
rect 8286 30796 8295 30856
rect 8985 30796 8994 30856
rect 9054 30796 9063 30856
rect 9753 30796 9762 30856
rect 9822 30796 9831 30856
rect 10521 30796 10530 30856
rect 10590 30796 10599 30856
rect 11289 30797 11298 30857
rect 11358 30797 11367 30857
rect 6690 30596 6750 30796
rect 7458 30596 7518 30796
rect 8226 30596 8286 30796
rect 8994 30596 9054 30796
rect 9762 30596 9822 30796
rect 10530 30596 10590 30796
rect 11298 30596 11358 30797
rect 12057 30796 12066 30856
rect 12126 30796 12135 30856
rect 12825 30796 12834 30856
rect 12894 30796 12903 30856
rect 13593 30796 13602 30856
rect 13662 30796 13671 30856
rect 14361 30796 14370 30856
rect 14430 30796 14439 30856
rect 15129 30796 15138 30856
rect 15198 30796 15207 30856
rect 15897 30796 15906 30856
rect 15966 30796 15975 30856
rect 16665 30796 16674 30856
rect 16734 30796 16743 30856
rect 17433 30796 17442 30856
rect 17502 30796 17511 30856
rect 18201 30796 18210 30856
rect 18270 30796 18279 30856
rect 18969 30796 18978 30856
rect 19038 30796 19047 30856
rect 19737 30796 19746 30856
rect 19806 30796 19815 30856
rect 20505 30796 20514 30856
rect 20574 30796 20583 30856
rect 21273 30796 21282 30856
rect 21342 30796 21351 30856
rect 22041 30796 22050 30856
rect 22110 30796 22119 30856
rect 22809 30796 22818 30856
rect 22878 30796 22887 30856
rect 23577 30796 23586 30856
rect 23646 30796 23655 30856
rect 30489 30796 30498 30856
rect 30558 30796 30567 30856
rect 31257 30797 31266 30857
rect 31326 30797 31335 30857
rect 12066 30596 12126 30796
rect 12834 30596 12894 30796
rect 13602 30596 13662 30796
rect 14370 30596 14430 30796
rect 15138 30596 15198 30796
rect 15906 30596 15966 30796
rect 16674 30596 16734 30796
rect 17442 30596 17502 30796
rect 18210 30596 18270 30796
rect 18978 30596 19038 30796
rect 19746 30596 19806 30796
rect 20514 30596 20574 30796
rect 21282 30596 21342 30796
rect 22050 30596 22110 30796
rect 22818 30596 22878 30796
rect 23586 30596 23646 30796
rect 24000 30596 24440 30605
rect 5922 30456 24000 30596
rect 24000 30447 24440 30456
rect 30498 30256 30558 30796
rect 30498 30187 30558 30196
rect 31266 29858 31326 30797
rect 32025 30796 32034 30856
rect 32094 30796 32103 30856
rect 32793 30796 32802 30856
rect 32862 30796 32871 30856
rect 33561 30796 33570 30856
rect 33630 30796 33639 30856
rect 34329 30796 34338 30856
rect 34398 30796 34407 30856
rect 35097 30796 35106 30856
rect 35166 30796 35175 30856
rect 35865 30796 35874 30856
rect 35934 30796 35943 30856
rect 31257 29798 31266 29858
rect 31326 29798 31335 29858
rect 31266 29797 31326 29798
rect 32034 29456 32094 30796
rect 32025 29396 32034 29456
rect 32094 29396 32103 29456
rect 32802 29056 32862 30796
rect 32793 28996 32802 29056
rect 32862 28996 32871 29056
rect 33570 28656 33630 30796
rect 33561 28596 33570 28656
rect 33630 28596 33639 28656
rect 34338 28256 34398 30796
rect 34329 28196 34338 28256
rect 34398 28196 34407 28256
rect 35106 27856 35166 30796
rect 35097 27796 35106 27856
rect 35166 27796 35175 27856
rect 35874 27456 35934 30796
rect 35865 27396 35874 27456
rect 35934 27396 35943 27456
rect 23991 26284 24000 26724
rect 24440 26284 24449 26724
rect 20 24776 200 24785
rect 200 24596 620 24776
rect 800 24596 809 24776
rect 20 24587 200 24596
<< via4 >>
rect 5922 30797 5982 30857
rect 6690 30796 6750 30856
rect 7458 30796 7518 30856
rect 8226 30796 8286 30856
rect 8994 30796 9054 30856
rect 9762 30796 9822 30856
rect 10530 30796 10590 30856
rect 11298 30797 11358 30857
rect 12066 30796 12126 30856
rect 12834 30796 12894 30856
rect 13602 30796 13662 30856
rect 14370 30796 14430 30856
rect 15138 30796 15198 30856
rect 15906 30796 15966 30856
rect 16674 30796 16734 30856
rect 17442 30796 17502 30856
rect 18210 30796 18270 30856
rect 18978 30796 19038 30856
rect 19746 30796 19806 30856
rect 20514 30796 20574 30856
rect 21282 30796 21342 30856
rect 22050 30796 22110 30856
rect 22818 30796 22878 30856
rect 23586 30796 23646 30856
rect 30498 30796 30558 30856
rect 31266 30797 31326 30857
rect 24000 30456 24440 30596
rect 32034 30796 32094 30856
rect 32802 30796 32862 30856
rect 33570 30796 33630 30856
rect 34338 30796 34398 30856
rect 35106 30796 35166 30856
rect 35874 30796 35934 30856
rect 24000 26284 24440 26724
rect 20 24596 200 24776
<< metal5 >>
rect 5922 30857 5982 30996
rect 5922 30788 5982 30797
rect 6690 30856 6750 30996
rect 6690 30787 6750 30796
rect 7458 30856 7518 30996
rect 7458 30787 7518 30796
rect 8226 30856 8286 30996
rect 8226 30787 8286 30796
rect 8994 30856 9054 30996
rect 8994 30787 9054 30796
rect 9762 30856 9822 30996
rect 9762 30787 9822 30796
rect 10530 30856 10590 30996
rect 10530 30787 10590 30796
rect 11298 30857 11358 30996
rect 11298 30788 11358 30797
rect 12066 30856 12126 30996
rect 12066 30787 12126 30796
rect 12834 30856 12894 30996
rect 12834 30787 12894 30796
rect 13602 30856 13662 30996
rect 13602 30787 13662 30796
rect 14370 30856 14430 30996
rect 14370 30787 14430 30796
rect 15138 30856 15198 30996
rect 15138 30787 15198 30796
rect 15906 30856 15966 30996
rect 15906 30787 15966 30796
rect 16674 30856 16734 30996
rect 16674 30787 16734 30796
rect 17442 30856 17502 30996
rect 17442 30787 17502 30796
rect 18210 30856 18270 30996
rect 18210 30787 18270 30796
rect 18978 30856 19038 30996
rect 18978 30787 19038 30796
rect 19746 30856 19806 30996
rect 19746 30787 19806 30796
rect 20514 30856 20574 30996
rect 20514 30787 20574 30796
rect 21282 30856 21342 30996
rect 21282 30787 21342 30796
rect 22050 30856 22110 30996
rect 22050 30787 22110 30796
rect 22818 30856 22878 30996
rect 22818 30787 22878 30796
rect 23586 30856 23646 30996
rect 24354 30796 24414 30996
rect 25122 30796 25182 30996
rect 25890 30796 25950 30996
rect 26658 30796 26718 30996
rect 27426 30796 27486 30996
rect 28194 30796 28254 30996
rect 28962 30796 29022 30996
rect 29730 30796 29790 30996
rect 30498 30856 30558 30996
rect 23586 30787 23646 30796
rect 30498 30787 30558 30796
rect 31266 30857 31326 30996
rect 31266 30788 31326 30797
rect 32034 30856 32094 30996
rect 32034 30787 32094 30796
rect 32802 30856 32862 30996
rect 32802 30787 32862 30796
rect 33570 30856 33630 30996
rect 33570 30787 33630 30796
rect 34338 30856 34398 30996
rect 34338 30787 34398 30796
rect 35106 30856 35166 30996
rect 35106 30787 35166 30796
rect 35874 30856 35934 30996
rect 36642 30796 36702 30996
rect 37410 30796 37470 30996
rect 38178 30796 38238 30996
rect 35874 30787 35934 30796
rect 23991 30456 24000 30596
rect 24440 30456 24449 30596
rect 24000 26724 24440 30456
rect 0 24596 20 24776
rect 200 24596 209 24776
rect 0 21396 200 21576
rect 0 18196 200 18376
rect 0 14996 200 15176
rect 24000 0 24440 26284
rect 24800 0 25240 30596
use r2r_dac  r2r_dac_0
timestamp 1746729020
transform -1 0 23462 0 -1 27417
box -89 -93 5515 1987
<< labels >>
flabel metal5 s 37410 30796 37470 30996 4 FreeSans 320 0 0 0 clk
port 2 nsew
flabel metal5 s 38178 30796 38238 30996 4 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal5 s 36642 30796 36702 30996 4 FreeSans 320 0 0 0 rst_n
port 4 nsew
flabel metal5 s 35874 30796 35934 30996 4 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew
flabel metal5 s 35106 30796 35166 30996 4 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew
flabel metal5 s 34338 30796 34398 30996 4 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew
flabel metal5 s 33570 30796 33630 30996 4 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew
flabel metal5 s 32802 30796 32862 30996 4 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew
flabel metal5 s 32034 30796 32094 30996 4 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew
flabel metal5 s 31266 30796 31326 30996 4 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew
flabel metal5 s 30498 30796 30558 30996 4 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew
flabel metal5 s 29730 30796 29790 30996 4 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew
flabel metal5 s 28962 30796 29022 30996 4 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew
flabel metal5 s 28194 30796 28254 30996 4 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew
flabel metal5 s 27426 30796 27486 30996 4 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew
flabel metal5 s 26658 30796 26718 30996 4 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew
flabel metal5 s 25890 30796 25950 30996 4 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew
flabel metal5 s 25122 30796 25182 30996 4 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew
flabel metal5 s 24354 30796 24414 30996 4 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew
flabel metal5 s 11298 30796 11358 30996 4 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew
flabel metal5 s 10530 30796 10590 30996 4 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew
flabel metal5 s 9762 30796 9822 30996 4 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew
flabel metal5 s 8994 30796 9054 30996 4 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew
flabel metal5 s 8226 30796 8286 30996 4 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew
flabel metal5 s 7458 30796 7518 30996 4 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew
flabel metal5 s 6690 30796 6750 30996 4 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew
flabel metal5 s 5922 30796 5982 30996 4 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew
flabel metal5 s 17442 30796 17502 30996 4 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew
flabel metal5 s 16674 30796 16734 30996 4 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew
flabel metal5 s 15906 30796 15966 30996 4 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew
flabel metal5 s 15138 30796 15198 30996 4 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew
flabel metal5 s 14370 30796 14430 30996 4 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew
flabel metal5 s 13602 30796 13662 30996 4 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew
flabel metal5 s 12834 30796 12894 30996 4 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew
flabel metal5 s 12066 30796 12126 30996 4 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew
flabel metal5 s 23586 30796 23646 30996 4 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew
flabel metal5 s 22818 30796 22878 30996 4 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew
flabel metal5 s 22050 30796 22110 30996 4 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew
flabel metal5 s 21282 30796 21342 30996 4 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew
flabel metal5 s 20514 30796 20574 30996 4 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew
flabel metal5 s 19746 30796 19806 30996 4 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew
flabel metal5 s 18978 30796 19038 30996 4 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew
flabel metal5 s 18210 30796 18270 30996 4 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew
flabel metal5 s 0 24596 200 24776 0 FreeSans 320 0 0 0 ua[0]
port 45 nsew
flabel metal5 s 0 21396 200 21576 0 FreeSans 320 0 0 0 ua[1]
port 46 nsew
flabel metal5 s 0 18196 200 18376 0 FreeSans 320 0 0 0 ua[2]
port 47 nsew
flabel metal5 s 0 14996 200 15176 0 FreeSans 320 0 0 0 ua[3]
port 48 nsew
flabel metal5 s 24000 0 24440 30596 0 FreeSans 320 0 0 0 VGND
port 49 nsew
flabel metal5 s 24800 0 25240 30596 0 FreeSans 320 0 0 0 VPWR
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 40416 30996
<< end >>
