magic
tech ihp-sg13g2
timestamp 1746820180
<< pwell >>
rect -1401 -512 1401 528
<< psubdiff >>
rect -1370 490 1370 497
rect -1370 474 -1324 490
rect 1324 474 1370 490
rect -1370 467 1370 474
rect -1370 451 -1340 467
rect -1370 -435 -1363 451
rect -1347 -435 -1340 451
rect -1370 -451 -1340 -435
rect 1340 451 1370 467
rect 1340 -435 1347 451
rect 1363 -435 1370 451
rect 1340 -451 1370 -435
rect -1370 -458 1370 -451
rect -1370 -474 -1324 -458
rect 1324 -474 1370 -458
rect -1370 -481 1370 -474
<< psubdiffcont >>
rect -1324 474 1324 490
rect -1363 -435 -1347 451
rect 1347 -435 1363 451
rect -1324 -474 1324 -458
<< metal1 >>
rect -1363 474 -1324 490
rect 1324 474 1363 490
rect -1363 451 -1347 474
rect -1363 -458 -1347 -435
rect 1347 451 1363 474
rect 1347 -458 1363 -435
rect -1363 -474 -1324 -458
rect 1324 -474 1363 -458
use rhigh  rhigh_0
timestamp 1746820100
transform 1 0 -1299 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_1
timestamp 1746820100
transform 1 0 -1201 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_2
timestamp 1746820100
transform 1 0 -1103 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_3
timestamp 1746820100
transform 1 0 -1005 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_4
timestamp 1746820100
transform 1 0 -907 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_5
timestamp 1746820100
transform 1 0 -809 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_6
timestamp 1746820100
transform 1 0 -711 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_7
timestamp 1746820100
transform 1 0 -613 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_8
timestamp 1746820100
transform 1 0 -515 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_9
timestamp 1746820100
transform 1 0 -417 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_10
timestamp 1746820100
transform 1 0 -319 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_11
timestamp 1746820100
transform 1 0 -221 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_12
timestamp 1746820100
transform 1 0 -123 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_13
timestamp 1746820100
transform 1 0 -25 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_14
timestamp 1746820100
transform 1 0 73 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_15
timestamp 1746820100
transform 1 0 171 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_16
timestamp 1746820100
transform 1 0 269 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_17
timestamp 1746820100
transform 1 0 367 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_18
timestamp 1746820100
transform 1 0 465 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_19
timestamp 1746820100
transform 1 0 563 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_20
timestamp 1746820100
transform 1 0 661 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_21
timestamp 1746820100
transform 1 0 759 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_22
timestamp 1746820100
transform 1 0 857 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_23
timestamp 1746820100
transform 1 0 955 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_24
timestamp 1746820100
transform 1 0 1053 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_25
timestamp 1746820100
transform 1 0 1151 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_26
timestamp 1746820100
transform 1 0 1249 0 1 -367
box 0 -43 50 793
<< labels >>
rlabel psubdiffcont 0 -466 0 -466 0 B
port 1 nsew
<< end >>
