magic
tech ihp-sg13g2
timestamp 1747416275
<< pwell >>
rect -1401 -512 1895 528
<< psubdiff >>
rect -1370 490 1864 497
rect -1370 474 -1324 490
rect 1818 474 1864 490
rect -1370 467 1864 474
rect -1370 451 -1340 467
rect -1370 -435 -1363 451
rect -1347 -435 -1340 451
rect -1370 -451 -1340 -435
rect 1834 451 1864 467
rect 1834 -435 1841 451
rect 1857 -435 1864 451
rect 1834 -451 1864 -435
rect -1370 -458 1864 -451
rect -1370 -474 -1324 -458
rect 1818 -474 1864 -458
rect -1370 -481 1864 -474
<< psubdiffcont >>
rect -1324 474 1818 490
rect -1363 -435 -1347 451
rect 1841 -435 1857 451
rect -1324 -474 1818 -458
<< metal1 >>
rect -1363 474 -1324 490
rect 1818 474 1857 490
rect -1363 451 -1347 474
rect -1363 -458 -1347 -435
rect 1841 451 1857 474
rect 1841 -458 1857 -435
rect -1363 -474 -1324 -458
rect 1818 -474 1857 -458
use rhigh  rhigh_0
timestamp 1746820100
transform 1 0 -1299 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_1
timestamp 1746820100
transform 1 0 -1182 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_2
timestamp 1746820100
transform 1 0 -1065 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_3
timestamp 1746820100
transform 1 0 -948 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_4
timestamp 1746820100
transform 1 0 -831 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_5
timestamp 1746820100
transform 1 0 -714 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_6
timestamp 1746820100
transform 1 0 -597 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_7
timestamp 1746820100
transform 1 0 -480 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_8
timestamp 1746820100
transform 1 0 -363 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_9
timestamp 1746820100
transform 1 0 -246 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_10
timestamp 1746820100
transform 1 0 -129 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_11
timestamp 1746820100
transform 1 0 -12 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_12
timestamp 1746820100
transform 1 0 105 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_13
timestamp 1746820100
transform 1 0 222 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_14
timestamp 1746820100
transform 1 0 339 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_15
timestamp 1746820100
transform 1 0 456 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_16
timestamp 1746820100
transform 1 0 573 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_17
timestamp 1746820100
transform 1 0 690 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_18
timestamp 1746820100
transform 1 0 807 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_19
timestamp 1746820100
transform 1 0 924 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_20
timestamp 1746820100
transform 1 0 1041 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_21
timestamp 1746820100
transform 1 0 1158 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_22
timestamp 1746820100
transform 1 0 1275 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_23
timestamp 1746820100
transform 1 0 1392 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_24
timestamp 1746820100
transform 1 0 1509 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_25
timestamp 1746820100
transform 1 0 1626 0 1 -367
box 0 -43 50 793
use rhigh  rhigh_26
timestamp 1746820100
transform 1 0 1743 0 1 -367
box 0 -43 50 793
<< labels >>
rlabel psubdiffcont 247 -466 247 -466 0 B
port 1 nsew
<< end >>
