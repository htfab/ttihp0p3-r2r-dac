magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747416626
<< metal1 >>
rect -13 197 215 1911
rect 349 1697 683 1783
rect 817 1697 1151 1784
rect 1285 1697 1619 1783
rect 1753 1697 1853 1783
rect 1519 1611 1619 1697
rect 1987 1611 2087 1783
rect 2221 1697 2555 1784
rect 2689 1697 3023 1783
rect 3157 1697 3257 1783
rect 1519 1525 2087 1611
rect 2923 1611 3023 1697
rect 3391 1611 3491 1783
rect 3625 1697 3959 1784
rect 4093 1697 4427 1783
rect 4561 1697 4661 1783
rect 2923 1525 3491 1611
rect 4327 1611 4427 1697
rect 4795 1611 4895 1783
rect 5029 1697 5363 1784
rect 5497 1697 5831 1783
rect 5965 1697 6065 1783
rect 4327 1525 4895 1611
rect 817 283 1385 369
rect 817 197 917 283
rect -13 111 449 197
rect 583 111 917 197
rect 1051 111 1151 197
rect 1285 111 1385 283
rect 2221 283 2789 369
rect 2221 197 2321 283
rect 1519 111 1853 197
rect 1987 111 2321 197
rect 2455 111 2555 197
rect 2689 111 2789 283
rect 3625 283 4193 369
rect 3625 197 3725 283
rect 2923 111 3257 197
rect 3391 111 3725 197
rect 3859 111 3959 197
rect 4093 111 4193 283
rect 5029 283 5597 369
rect 5029 197 5129 283
rect 4327 111 4661 197
rect 4795 111 5129 197
rect 5263 111 5363 197
rect 5497 111 5597 283
rect 5731 111 6065 197
rect -13 -17 215 111
rect 6199 -17 6427 1911
use resistors  resistors_0
timestamp 1747416275
transform 1 0 2713 0 1 931
box -2802 -1024 3790 1056
<< labels >>
flabel metal1 349 111 449 197 0 FreeSans 256 0 0 0 GND
port 1 nsew ground bidirectional
flabel metal1 1051 111 1151 197 0 FreeSans 256 0 0 0 IN[0]
port 2 nsew signal input
flabel metal1 1753 1697 1853 1783 0 FreeSans 256 0 0 0 IN[1]
port 3 nsew signal input
flabel metal1 2455 111 2555 197 0 FreeSans 256 0 0 0 IN[2]
port 4 nsew signal input
flabel metal1 3157 1697 3257 1783 0 FreeSans 256 0 0 0 IN[3]
port 5 nsew signal input
flabel metal1 3859 111 3959 197 0 FreeSans 256 0 0 0 IN[4]
port 6 nsew signal input
flabel metal1 4561 1697 4661 1783 0 FreeSans 256 0 0 0 IN[5]
port 7 nsew signal input
flabel metal1 5263 111 5363 197 0 FreeSans 256 0 0 0 IN[6]
port 8 nsew signal input
flabel metal1 5965 1697 6065 1783 0 FreeSans 256 0 0 0 IN[7]
port 9 nsew signal input
flabel metal1 5497 1697 5831 1783 0 FreeSans 256 0 0 0 OUT
port 10 nsew signal output
<< end >>
