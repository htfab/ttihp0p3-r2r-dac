magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747591589
<< metal1 >>
rect -48 197 215 1946
rect 362 1697 709 1783
rect 856 1697 1203 1784
rect 1350 1697 1697 1783
rect 1844 1697 1944 1783
rect 1597 1611 1697 1697
rect 2091 1611 2191 1783
rect 2338 1697 2685 1784
rect 2832 1697 3179 1783
rect 3326 1697 3426 1783
rect 1597 1525 2191 1611
rect 3079 1611 3179 1697
rect 3573 1611 3673 1783
rect 3820 1697 4167 1784
rect 4314 1697 4661 1783
rect 4808 1697 4908 1783
rect 3079 1525 3673 1611
rect 4561 1611 4661 1697
rect 5055 1611 5155 1783
rect 5302 1697 5649 1784
rect 5796 1697 6143 1783
rect 6290 1697 6390 1783
rect 4561 1525 5155 1611
rect 856 283 1450 369
rect 856 197 956 283
rect -48 111 462 197
rect 609 111 956 197
rect 1103 111 1203 197
rect 1350 111 1450 283
rect 2338 283 2932 369
rect 2338 197 2438 283
rect 1597 111 1944 197
rect 2091 111 2438 197
rect 2585 111 2685 197
rect 2832 111 2932 283
rect 3820 283 4414 369
rect 3820 197 3920 283
rect 3079 111 3426 197
rect 3573 111 3920 197
rect 4067 111 4167 197
rect 4314 111 4414 283
rect 5302 283 5896 369
rect 5302 197 5402 283
rect 4561 111 4908 197
rect 5055 111 5402 197
rect 5549 111 5649 197
rect 5796 111 5896 283
rect 6043 111 6390 197
rect -48 -52 215 111
rect 6537 -52 6800 1946
use resistors  resistors_0
timestamp 1747591324
transform 1 0 2713 0 1 931
box -2837 -1059 4163 1091
<< labels >>
flabel metal1 362 111 462 197 0 FreeSans 256 0 0 0 GND
port 1 nsew ground bidirectional
flabel metal1 1103 111 1203 197 0 FreeSans 256 0 0 0 IN[0]
port 2 nsew signal input
flabel metal1 1844 1697 1944 1783 0 FreeSans 256 0 0 0 IN[1]
port 3 nsew signal input
flabel metal1 2585 111 2685 197 0 FreeSans 256 0 0 0 IN[2]
port 4 nsew signal input
flabel metal1 3326 1697 3426 1783 0 FreeSans 256 0 0 0 IN[3]
port 5 nsew signal input
flabel metal1 4067 111 4167 197 0 FreeSans 256 0 0 0 IN[4]
port 6 nsew signal input
flabel metal1 4808 1697 4908 1783 0 FreeSans 256 0 0 0 IN[5]
port 7 nsew signal input
flabel metal1 5549 111 5649 197 0 FreeSans 256 0 0 0 IN[6]
port 8 nsew signal input
flabel metal1 5796 1697 6143 1783 0 FreeSans 256 0 0 0 OUT
port 10 nsew signal output
flabel metal1 6290 1697 6390 1783 0 FreeSans 256 0 0 0 IN[7]
port 9 nsew signal input
<< end >>
