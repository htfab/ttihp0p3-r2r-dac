magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747591324
<< pwell >>
rect -2837 -1059 4163 1091
<< psubdiff >>
rect -2775 1015 4101 1029
rect -2775 983 -2683 1015
rect 4009 983 4101 1015
rect -2775 969 4101 983
rect -2775 937 -2715 969
rect -2775 -905 -2761 937
rect -2729 -905 -2715 937
rect -2775 -937 -2715 -905
rect 4041 937 4101 969
rect 4041 -905 4055 937
rect 4087 -905 4101 937
rect 4041 -937 4101 -905
rect -2775 -951 4101 -937
rect -2775 -983 -2683 -951
rect 4009 -983 4101 -951
rect -2775 -997 4101 -983
<< psubdiffcont >>
rect -2683 983 4009 1015
rect -2761 -905 -2729 937
rect 4055 -905 4087 937
rect -2683 -983 4009 -951
<< metal1 >>
rect -2761 983 -2683 1015
rect 4009 983 4087 1015
rect -2761 937 -2729 983
rect -2761 -951 -2729 -905
rect 4055 937 4087 983
rect 4055 -951 4087 -905
rect -2761 -983 -2683 -951
rect 4009 -983 4087 -951
use rhigh  rhigh_0
timestamp 1746820100
transform 1 0 -2598 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_1
timestamp 1746820100
transform 1 0 -2351 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_2
timestamp 1746820100
transform 1 0 -2104 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_3
timestamp 1746820100
transform 1 0 -1857 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_4
timestamp 1746820100
transform 1 0 -1610 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_5
timestamp 1746820100
transform 1 0 -1363 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_6
timestamp 1746820100
transform 1 0 -1116 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_7
timestamp 1746820100
transform 1 0 -869 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_8
timestamp 1746820100
transform 1 0 -622 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_9
timestamp 1746820100
transform 1 0 -375 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_10
timestamp 1746820100
transform 1 0 -128 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_11
timestamp 1746820100
transform 1 0 119 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_12
timestamp 1746820100
transform 1 0 366 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_13
timestamp 1746820100
transform 1 0 613 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_14
timestamp 1746820100
transform 1 0 860 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_15
timestamp 1746820100
transform 1 0 1107 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_16
timestamp 1746820100
transform 1 0 1354 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_17
timestamp 1746820100
transform 1 0 1601 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_18
timestamp 1746820100
transform 1 0 1848 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_19
timestamp 1746820100
transform 1 0 2095 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_20
timestamp 1746820100
transform 1 0 2342 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_21
timestamp 1746820100
transform 1 0 2589 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_22
timestamp 1746820100
transform 1 0 2836 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_23
timestamp 1746820100
transform 1 0 3083 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_24
timestamp 1746820100
transform 1 0 3330 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_25
timestamp 1746820100
transform 1 0 3577 0 1 -734
box 0 -86 100 1586
use rhigh  rhigh_26
timestamp 1746820100
transform 1 0 3824 0 1 -734
box 0 -86 100 1586
<< labels >>
rlabel psubdiffcont 663 -967 663 -967 0 B
port 1 nsew
<< end >>
